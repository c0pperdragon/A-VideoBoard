package VICTypes is    -- untested...

   type t_VICType is (CLOCKS63, CLOCKS64, CLOCKS65);

end VICTypes;
